module tweakablecipher (/*AUTOARG*/ ) ;
   output [63+64*fullcnt:0] nextcnt;
   output [127:0] 	       nextkey, nexttweak, nextstate;
   
endmodule // tweakablecipher
