module padding_decider (/*AUTOARG*/ ) ;
`include "romulus_config_pkg.v"

   input  [15:0] fsm;
   input [CNTW-1:0] cnt;
   input [15:0]     seglen;

   generate begin
      if (ز)
      if (TBC == DUMMY) begin
         always @ (*) begin
            
         end
      end
   end

endmodule // padding_decider

